process(a,b)
begin
 if (a <> b) then
 c <= '0';
 else
 c <= '1';
 end if;
end process;